library IEEE;
use IEEE.std_logic_1164.all;
use work.HermesPackage.all;

entity testbench is
	generic(
		X_NODES: integer := 1;
		Y_NODES: integer := 1
	);
end entity;

architecture behavioral of testbench is
	signal clock: std_logic := '0';
	signal reset: std_logic;

	signal clock_tx:	regNport;
	signal tx:			regNport;
	signal data_out:	arrayNport_regflit;
	signal credit_i:	regNport;

	signal credit_o:	regNport;
	signal rx:			regNport;

	constant NB_ROUTERS : integer :=  X_NODES * Y_NODES;

	signal data_in:	array_buffer;
	signal data_ack:	port_buffer;
	signal data_av:		port_buffer;

-----------------------------------------------------------------

	signal address1, data1: std_logic_vector(15 downto 0);
	signal ce1: std_logic;

	type packet is array (0 to 16) of std_logic_vector(15 downto 0);
	constant pck1 : packet := 
	(
		x"0000", x"000F", x"1001", x"2002", x"3003", x"4004", x"5005",
		x"6006", x"7007", x"8008", x"9009", x"A00A",
		x"B00B", x"C00C", x"D00D", x"E00E", x"F00F"
	);
begin
	reset <= '1', '0' after 15 ns;
	clock <= not clock after 10 ns;

	cu: for i in 0 to NPORT - 1 generate
		clock_tx(i) <= clock;
	end generate;

	node1:	entity	work.node
	port map(
		clock => clock,
		reset => reset,

		clock_rx => clock_tx,
		rx =>	tx,
		data_in => data_out,
		credit_o => credit_i,

		data_out => data_in,
		data_ack => data_ack,
		data_av => data_av
	);

	--------------------


	process(reset, clock)
	begin
		if reset='1' then
			tx <= (others => '0');
		elsif rising_edge(clock) then
			if ce1='1' and address1=x"FFFF" then
				tx(LOCAL) <= '1';
				data_out(LOCAL) <= data1;

			elsif credit_i(LOCAL) = '1' then -- important: flow control
				tx(LOCAL) <= '0';
			end if;
		end if;
	end process;

	address1 <= x"FFFF"; -- address generated by the processor
	process
		variable i : integer:= 0;
	begin
		ce1 <= '0';
		wait for 400 ns; -- time between packets
		i := 0;
		while i < 17 loop
			if credit_i(LOCAL) = '1' then -- important: flow control
				data1 <= pck1(i); -- simulate a write( pck(i), address_noc)
				ce1 <= '1';
				wait for 20 ns;
				ce1 <= '0';
				wait for 20 ns;
				i := i + 1;
			else
				wait for 20 ns;
			end if;
		end loop;
	end process;


end architecture;